//interfaces
`include "interface.svh"

//package
`include "packages.sv"

//rtl
`include "without_pipelining.sv"
`include "pipelined_without_forwarding.sv"
`include "pipelined_with_forwarding.sv"
`include "top.sv"